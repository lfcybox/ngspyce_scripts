**.subckt nmos_tb
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
**** begin user architecture code

.temp 27
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice ss
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice ff
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice sf
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice fs



Vg G 0 1.8
Vs S 0 0
Vd D 0 1.8
Vb B 0 0

.save v(G) v(D) v(S) v(B)
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gmbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vgs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[css]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbs]


**** end user architecture code
**.ends
** flattened .save nodes
.save v(G) v(D) v(S) v(B)
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gmbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vgs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[css]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[csb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cbb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbs]
.end
