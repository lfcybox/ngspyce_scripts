* bjt corner test http://ngspice.sourceforge.net/ngspice-tutorial.html
* Using UPPERCASE labels such as SIM_TEMP and SIM_BJTCORNER
* as placeholders for ngspyce to replace to sweep corners,
* temperature, etc.

*.lib corner_test.lib typ
*.lib corner_test.lib betalow

.lib corner_test.lib SIM_BJTCORNER
*.temp SIM_TEMP

R3 vcc intc 10k
R1 vcc intb 68k
R2 intb 0 10k
Cout out intc 10u
Cin intb in 10u
VCC vcc 0 5
Vin in 0 dc 0 ac 1 sin(0 1m 500)
RLoad out 0 100k
Q1 intc intb 0 BC546B

*.tran 10u 10m

.end
