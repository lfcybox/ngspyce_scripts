**.subckt test_sch2
R1 OUT IN1 100k m=1
R2 IN2 OUT 50k m=1
V1 IN1 GND 3
V2 IN2 GND 3
**.ends
.GLOBAL GND
** flattened .save nodes
.end
