**.subckt test_sky_rc
XC1 OUT GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=2 m=2
V1 IN GND pulse 0 3 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 ' 
XR2 GND OUT GND sky130_fd_pr__res_xhigh_po W=1 L=1000 mult=1 m=1
XR3 OUT IN GND sky130_fd_pr__res_xhigh_po W=1 L=1000 mult=1 m=1
**** begin user architecture code

.temp 27
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice ss
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice ff
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice sf
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice fs

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
